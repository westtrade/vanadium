module utils

units := ["h", "m", "s", "ms", "μs", "ns"]
divisors := [3_600_000.0, 60_000.0, 1_000.0, 1.0, 1e-3, 1e-6]
